----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:59:36 12/12/2020 
-- Design Name: 
-- Module Name:    CharacterIn7Seg - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CharacterIn7Seg is
	port(
		sel: in std_logic_vector(1 downto 0);
		segment_out: out std_logic_vector(7 downto 0)
	);
end CharacterIn7Seg;

architecture Behavioral of CharacterIn7Seg is

begin
	with sel select segment_out <=
		"11101110" when "00",
		"00111110" when "01",
		"00011010" when "10",
		"01111010" when "11";

end Behavioral;

